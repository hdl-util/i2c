module master_tb ();
endmodule

